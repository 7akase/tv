`timescale 1ns / 1ps

`define ms *(1000`us)
`define us *(1000`ns)
`define ns *(1)
